// Copyright 2018 ETH Zurich and University of Bologna.
// Copyright and related rights are licensed under the Solderpad Hardware
// License, Version 0.51 (the "License"); you may not use this file except in
// compliance with the License.  You may obtain a copy of the License at
// http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
// or agreed to in writing, software, hardware and materials distributed under
// this License is distributed on an "AS IS" BASIS, WITHOUT WARRANTIES OR
// CONDITIONS OF ANY KIND, either express or implied. See the License for the
// specific language governing permissions and limitations under the License.

////////////////////////////////////////////////////////////////////////////////
//                                                                            //
// Authors:        Renzo Andri - andrire@student.ethz.ch                      //
//                 Igor Loi - igor.loi@unibo.it                               //
//                 Andreas Traber - atraber@student.ethz.ch                   //
//                 Sven Stucki - svstucki@student.ethz.ch                     //
//                 Michael Gautschi - gautschi@iis.ee.ethz.ch                 //
//                 Davide Schiavone - pschiavo@iis.ee.ethz.ch                 //
//                 Halfdan Bechmann - halfdan.bechmann@silabs.com             //
//                                                                            //
// Description:    RTL assertions for the id_stage module                     //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////


module cv32e40x_id_stage_sva
  import uvm_pkg::*;
  import cv32e40x_pkg::*;
(
  input logic           clk,
  input logic           rst_n,

  input logic [31:0]    instr,
  input logic           rf_we,
  input logic           alu_en,
  input logic           mul_en,
  input logic           lsu_en,
  input logic           wfi_insn,
  input logic           ebrk_insn,
  input logic           mret_insn,
  input logic           dret_insn,
  input logic           ecall_insn,
  input logic           fencei_insn,
  input logic           ex_ready_i,
  input logic           illegal_insn,
  input csr_opcode_e    csr_op,
  input if_id_pipe_t    if_id_pipe_i,
  input id_ex_pipe_t    id_ex_pipe_o,
  input logic           id_ready_o,
  input logic           id_valid_o,
  input ctrl_fsm_t      ctrl_fsm_i,
  input logic           xif_insn_accept,
  input logic [1:0]     rf_re
);


    // the instruction delivered to the ID stage should always be valid
    a_valid_instr :
      assert property (@(posedge clk)
                       (if_id_pipe_i.instr_valid & (~if_id_pipe_i.illegal_c_insn)) |-> (!$isunknown(instr)) )
        else `uvm_error("id_stage", $sformatf("%t, Instruction is valid, but has at least one X", $time));
/* todo: check and fix/remove
      // Check that instruction after taken branch is flushed (more should actually be flushed, but that is not checked here)
      // and that EX stage is ready to receive flushed instruction immediately
      property p_branch_taken_ex;
        @(posedge clk) disable iff (!rst_n) (branch_taken_ex == 1'b1) |-> ((ex_ready_i == 1'b1) &&
                                                                           (alu_en == 1'b0) &&
                                                                           (mul_en == 1'b0) &&
                                                                           (rf_we == 1'b0) &&
                                                                           (lsu_en == 1'b0));
      endproperty

      a_branch_taken_ex : assert property(p_branch_taken_ex) else `uvm_error("id_stage", "Assertion p_branch_taken_ex failed")
*/

/* todo: check and fix/remove
      // Check that if IRQ PC update does not coincide with IRQ related CSR write
      // MIE is excluded from the check because it has a bypass.
      property p_irq_csr;
        @(posedge clk) disable iff (!rst_n)
          (pc_set_o && (pc_mux_o == PC_EXCEPTION) &&
           ((exc_pc_mux_o == EXC_PC_EXCEPTION) || (exc_pc_mux_o == EXC_PC_IRQ)) &&
           id_ex_pipe_o.csr_access && (id_ex_pipe_o.csr_op != CSR_OP_READ)) |->
                                  ((id_ex_pipe_o.alu_operand_b[11:0] != CSR_MSTATUS) &&
                                   (id_ex_pipe_o.alu_operand_b[11:0] != CSR_MEPC) &&
                                   (id_ex_pipe_o.alu_operand_b[11:0] != CSR_MCAUSE) &&
                                   (id_ex_pipe_o.alu_operand_b[11:0] != CSR_MTVEC));
      endproperty

      a_irq_csr : assert property(p_irq_csr) else `uvm_error("id_stage", "Assertion p_irq_csr failed")
*/

/* todo: fix
      generate
        if (!A_EXTENSION) begin : gen_no_a_extension_assertions

          // Check that A extension opcodes are decoded as illegal when A extension not enabled
          property p_illegal_0;
          @(posedge clk) disable iff (!rst_n) (instr[6:0] == OPCODE_AMO) |-> (illegal_insn == 'b1);
        endproperty

          a_illegal_0 : assert property(p_illegal_0) else `uvm_error("id_stage", "Assertion p_illegal_0 failed")

        end
      endgenerate
*/
      // Check that illegal instruction has no other side effects
      // If xif accepts instruction, rf_we may still be 1
      property p_illegal_2;
        @(posedge clk) disable iff (!rst_n) (illegal_insn == 1'b1) |-> !(ebrk_insn || mret_insn || dret_insn ||
                                                                         ecall_insn || wfi_insn || fencei_insn ||
                                                                         alu_en || mul_en ||
                                                                         (rf_we && !xif_insn_accept) ||
                                                                         csr_op != CSR_OP_READ || lsu_en);
      endproperty

      a_illegal_2 : assert property(p_illegal_2) else `uvm_error("id_stage", "Assertion p_illegal_2 failed")

  // Halt implies not ready and not valid
  a_halt :
    assert property (@(posedge clk) disable iff (!rst_n)
                      (ctrl_fsm_i.halt_id && !ctrl_fsm_i.kill_id)
                      |-> (!id_ready_o && !id_valid_o))
      else `uvm_error("id_stage", "Halt should imply not ready and not valid")

  // Kill implies ready and not valid
  a_kill :
    assert property (@(posedge clk) disable iff (!rst_n)
                      (ctrl_fsm_i.kill_id)
                      |-> (id_ready_o && !id_valid_o))
      else `uvm_error("id_stage", "Kill should imply ready and not valid")
  
  // TODO: These may not be 100% correct in case
  // some instr bits are not clocked, and illegal insn would not be detected for example
  //   Could use full decoder in sva, and give it ungated instruction words
  // If decoder sets rf_re[0], if_id_pipe_i.rs1_enable must also be set
  a_predecoded_rf_re_0 :
  assert property (@(posedge clk) disable iff (!rst_n)
                    (rf_re[0] && if_id_pipe_i.instr_valid |-> if_id_pipe_i.rs1_enable))
    else `uvm_error("id_stage", "Predecoded rf_re[0] does not match decoder rf_re[0]")

  // If decoder sets rf_re[0], if_id_pipe_i.rs1_enable must also be set
  a_predecoded_rf_re_1 :
  assert property (@(posedge clk) disable iff (!rst_n)
                    (rf_re[1] && if_id_pipe_i.instr_valid |-> if_id_pipe_i.rs2_enable))
    else `uvm_error("id_stage", "Predecoded rf_re[0] does not match decoder rf_re[0]")
  
  // Illegal instruction must read all operands
  a_illegal_rs_enable:
  assert property (@(posedge clk) disable iff (!rst_n)
                    illegal_insn |->
                    (if_id_pipe_i.rs1_enable && if_id_pipe_i.rs2_enable))
    else `uvm_error ("id_stage", "Operands not enabled for illegal instruction")

  // rs2_enable can only be 1 if rs1_enable is also 1
  a_rs2_and_rs1 :
  assert property (@(posedge clk) disable iff (!rst_n)
                    (if_id_pipe_i.rs2_enable |-> if_id_pipe_i.rs1_enable))
    else `uvm_error("id_stage", "rs2_enable == 1 while rs1_enable == 0")


endmodule // cv32e40x_id_stage_sva

